module sinTable(input clk, input [9:0] addr, output reg [15:0] data);
reg [15:0] mem [0:1023];
initial mem[0] = 16'h0;
initial mem[1] = 16'hc9;
initial mem[2] = 16'h192;
initial mem[3] = 16'h25b;
initial mem[4] = 16'h324;
initial mem[5] = 16'h3ed;
initial mem[6] = 16'h4b6;
initial mem[7] = 16'h57e;
initial mem[8] = 16'h647;
initial mem[9] = 16'h710;
initial mem[10] = 16'h7d9;
initial mem[11] = 16'h8a1;
initial mem[12] = 16'h96a;
initial mem[13] = 16'ha32;
initial mem[14] = 16'hafb;
initial mem[15] = 16'hbc3;
initial mem[16] = 16'hc8b;
initial mem[17] = 16'hd53;
initial mem[18] = 16'he1b;
initial mem[19] = 16'hee3;
initial mem[20] = 16'hfab;
initial mem[21] = 16'h1072;
initial mem[22] = 16'h1139;
initial mem[23] = 16'h1200;
initial mem[24] = 16'h12c7;
initial mem[25] = 16'h138e;
initial mem[26] = 16'h1455;
initial mem[27] = 16'h151b;
initial mem[28] = 16'h15e1;
initial mem[29] = 16'h16a7;
initial mem[30] = 16'h176d;
initial mem[31] = 16'h1833;
initial mem[32] = 16'h18f8;
initial mem[33] = 16'h19bd;
initial mem[34] = 16'h1a82;
initial mem[35] = 16'h1b46;
initial mem[36] = 16'h1c0b;
initial mem[37] = 16'h1ccf;
initial mem[38] = 16'h1d93;
initial mem[39] = 16'h1e56;
initial mem[40] = 16'h1f19;
initial mem[41] = 16'h1fdc;
initial mem[42] = 16'h209f;
initial mem[43] = 16'h2161;
initial mem[44] = 16'h2223;
initial mem[45] = 16'h22e4;
initial mem[46] = 16'h23a6;
initial mem[47] = 16'h2467;
initial mem[48] = 16'h2527;
initial mem[49] = 16'h25e7;
initial mem[50] = 16'h26a7;
initial mem[51] = 16'h2767;
initial mem[52] = 16'h2826;
initial mem[53] = 16'h28e5;
initial mem[54] = 16'h29a3;
initial mem[55] = 16'h2a61;
initial mem[56] = 16'h2b1e;
initial mem[57] = 16'h2bdb;
initial mem[58] = 16'h2c98;
initial mem[59] = 16'h2d54;
initial mem[60] = 16'h2e10;
initial mem[61] = 16'h2ecc;
initial mem[62] = 16'h2f86;
initial mem[63] = 16'h3041;
initial mem[64] = 16'h30fb;
initial mem[65] = 16'h31b4;
initial mem[66] = 16'h326d;
initial mem[67] = 16'h3326;
initial mem[68] = 16'h33de;
initial mem[69] = 16'h3496;
initial mem[70] = 16'h354d;
initial mem[71] = 16'h3603;
initial mem[72] = 16'h36b9;
initial mem[73] = 16'h376f;
initial mem[74] = 16'h3824;
initial mem[75] = 16'h38d8;
initial mem[76] = 16'h398c;
initial mem[77] = 16'h3a3f;
initial mem[78] = 16'h3af2;
initial mem[79] = 16'h3ba4;
initial mem[80] = 16'h3c56;
initial mem[81] = 16'h3d07;
initial mem[82] = 16'h3db7;
initial mem[83] = 16'h3e67;
initial mem[84] = 16'h3f16;
initial mem[85] = 16'h3fc5;
initial mem[86] = 16'h4073;
initial mem[87] = 16'h4120;
initial mem[88] = 16'h41cd;
initial mem[89] = 16'h4279;
initial mem[90] = 16'h4325;
initial mem[91] = 16'h43d0;
initial mem[92] = 16'h447a;
initial mem[93] = 16'h4523;
initial mem[94] = 16'h45cc;
initial mem[95] = 16'h4674;
initial mem[96] = 16'h471c;
initial mem[97] = 16'h47c3;
initial mem[98] = 16'h4869;
initial mem[99] = 16'h490e;
initial mem[100] = 16'h49b3;
initial mem[101] = 16'h4a57;
initial mem[102] = 16'h4afa;
initial mem[103] = 16'h4b9d;
initial mem[104] = 16'h4c3f;
initial mem[105] = 16'h4ce0;
initial mem[106] = 16'h4d80;
initial mem[107] = 16'h4e20;
initial mem[108] = 16'h4ebf;
initial mem[109] = 16'h4f5d;
initial mem[110] = 16'h4ffa;
initial mem[111] = 16'h5097;
initial mem[112] = 16'h5133;
initial mem[113] = 16'h51ce;
initial mem[114] = 16'h5268;
initial mem[115] = 16'h5301;
initial mem[116] = 16'h539a;
initial mem[117] = 16'h5432;
initial mem[118] = 16'h54c9;
initial mem[119] = 16'h555f;
initial mem[120] = 16'h55f4;
initial mem[121] = 16'h5689;
initial mem[122] = 16'h571d;
initial mem[123] = 16'h57b0;
initial mem[124] = 16'h5842;
initial mem[125] = 16'h58d3;
initial mem[126] = 16'h5963;
initial mem[127] = 16'h59f3;
initial mem[128] = 16'h5a81;
initial mem[129] = 16'h5b0f;
initial mem[130] = 16'h5b9c;
initial mem[131] = 16'h5c28;
initial mem[132] = 16'h5cb3;
initial mem[133] = 16'h5d3d;
initial mem[134] = 16'h5dc6;
initial mem[135] = 16'h5e4f;
initial mem[136] = 16'h5ed6;
initial mem[137] = 16'h5f5d;
initial mem[138] = 16'h5fe2;
initial mem[139] = 16'h6067;
initial mem[140] = 16'h60eb;
initial mem[141] = 16'h616e;
initial mem[142] = 16'h61f0;
initial mem[143] = 16'h6271;
initial mem[144] = 16'h62f1;
initial mem[145] = 16'h6370;
initial mem[146] = 16'h63ee;
initial mem[147] = 16'h646b;
initial mem[148] = 16'h64e7;
initial mem[149] = 16'h6562;
initial mem[150] = 16'h65dd;
initial mem[151] = 16'h6656;
initial mem[152] = 16'h66ce;
initial mem[153] = 16'h6745;
initial mem[154] = 16'h67bc;
initial mem[155] = 16'h6831;
initial mem[156] = 16'h68a5;
initial mem[157] = 16'h6919;
initial mem[158] = 16'h698b;
initial mem[159] = 16'h69fc;
initial mem[160] = 16'h6a6c;
initial mem[161] = 16'h6adb;
initial mem[162] = 16'h6b4a;
initial mem[163] = 16'h6bb7;
initial mem[164] = 16'h6c23;
initial mem[165] = 16'h6c8e;
initial mem[166] = 16'h6cf8;
initial mem[167] = 16'h6d61;
initial mem[168] = 16'h6dc9;
initial mem[169] = 16'h6e30;
initial mem[170] = 16'h6e95;
initial mem[171] = 16'h6efa;
initial mem[172] = 16'h6f5e;
initial mem[173] = 16'h6fc0;
initial mem[174] = 16'h7022;
initial mem[175] = 16'h7082;
initial mem[176] = 16'h70e1;
initial mem[177] = 16'h7140;
initial mem[178] = 16'h719d;
initial mem[179] = 16'h71f9;
initial mem[180] = 16'h7254;
initial mem[181] = 16'h72ae;
initial mem[182] = 16'h7306;
initial mem[183] = 16'h735e;
initial mem[184] = 16'h73b5;
initial mem[185] = 16'h740a;
initial mem[186] = 16'h745e;
initial mem[187] = 16'h74b1;
initial mem[188] = 16'h7503;
initial mem[189] = 16'h7554;
initial mem[190] = 16'h75a4;
initial mem[191] = 16'h75f3;
initial mem[192] = 16'h7640;
initial mem[193] = 16'h768d;
initial mem[194] = 16'h76d8;
initial mem[195] = 16'h7722;
initial mem[196] = 16'h776b;
initial mem[197] = 16'h77b3;
initial mem[198] = 16'h77f9;
initial mem[199] = 16'h783f;
initial mem[200] = 16'h7883;
initial mem[201] = 16'h78c6;
initial mem[202] = 16'h7908;
initial mem[203] = 16'h7949;
initial mem[204] = 16'h7989;
initial mem[205] = 16'h79c7;
initial mem[206] = 16'h7a04;
initial mem[207] = 16'h7a41;
initial mem[208] = 16'h7a7c;
initial mem[209] = 16'h7ab5;
initial mem[210] = 16'h7aee;
initial mem[211] = 16'h7b25;
initial mem[212] = 16'h7b5c;
initial mem[213] = 16'h7b91;
initial mem[214] = 16'h7bc4;
initial mem[215] = 16'h7bf7;
initial mem[216] = 16'h7c29;
initial mem[217] = 16'h7c59;
initial mem[218] = 16'h7c88;
initial mem[219] = 16'h7cb6;
initial mem[220] = 16'h7ce2;
initial mem[221] = 16'h7d0e;
initial mem[222] = 16'h7d38;
initial mem[223] = 16'h7d61;
initial mem[224] = 16'h7d89;
initial mem[225] = 16'h7db0;
initial mem[226] = 16'h7dd5;
initial mem[227] = 16'h7df9;
initial mem[228] = 16'h7e1c;
initial mem[229] = 16'h7e3e;
initial mem[230] = 16'h7e5e;
initial mem[231] = 16'h7e7e;
initial mem[232] = 16'h7e9c;
initial mem[233] = 16'h7eb9;
initial mem[234] = 16'h7ed4;
initial mem[235] = 16'h7eef;
initial mem[236] = 16'h7f08;
initial mem[237] = 16'h7f20;
initial mem[238] = 16'h7f37;
initial mem[239] = 16'h7f4c;
initial mem[240] = 16'h7f61;
initial mem[241] = 16'h7f74;
initial mem[242] = 16'h7f86;
initial mem[243] = 16'h7f96;
initial mem[244] = 16'h7fa6;
initial mem[245] = 16'h7fb4;
initial mem[246] = 16'h7fc1;
initial mem[247] = 16'h7fcd;
initial mem[248] = 16'h7fd7;
initial mem[249] = 16'h7fe0;
initial mem[250] = 16'h7fe8;
initial mem[251] = 16'h7fef;
initial mem[252] = 16'h7ff5;
initial mem[253] = 16'h7ff9;
initial mem[254] = 16'h7ffc;
initial mem[255] = 16'h7ffe;
initial mem[256] = 16'h7fff;
initial mem[257] = 16'h7ffe;
initial mem[258] = 16'h7ffc;
initial mem[259] = 16'h7ff9;
initial mem[260] = 16'h7ff5;
initial mem[261] = 16'h7fef;
initial mem[262] = 16'h7fe8;
initial mem[263] = 16'h7fe0;
initial mem[264] = 16'h7fd7;
initial mem[265] = 16'h7fcd;
initial mem[266] = 16'h7fc1;
initial mem[267] = 16'h7fb4;
initial mem[268] = 16'h7fa6;
initial mem[269] = 16'h7f96;
initial mem[270] = 16'h7f86;
initial mem[271] = 16'h7f74;
initial mem[272] = 16'h7f61;
initial mem[273] = 16'h7f4c;
initial mem[274] = 16'h7f37;
initial mem[275] = 16'h7f20;
initial mem[276] = 16'h7f08;
initial mem[277] = 16'h7eef;
initial mem[278] = 16'h7ed4;
initial mem[279] = 16'h7eb9;
initial mem[280] = 16'h7e9c;
initial mem[281] = 16'h7e7e;
initial mem[282] = 16'h7e5e;
initial mem[283] = 16'h7e3e;
initial mem[284] = 16'h7e1c;
initial mem[285] = 16'h7df9;
initial mem[286] = 16'h7dd5;
initial mem[287] = 16'h7db0;
initial mem[288] = 16'h7d89;
initial mem[289] = 16'h7d61;
initial mem[290] = 16'h7d38;
initial mem[291] = 16'h7d0e;
initial mem[292] = 16'h7ce2;
initial mem[293] = 16'h7cb6;
initial mem[294] = 16'h7c88;
initial mem[295] = 16'h7c59;
initial mem[296] = 16'h7c29;
initial mem[297] = 16'h7bf7;
initial mem[298] = 16'h7bc4;
initial mem[299] = 16'h7b91;
initial mem[300] = 16'h7b5c;
initial mem[301] = 16'h7b25;
initial mem[302] = 16'h7aee;
initial mem[303] = 16'h7ab5;
initial mem[304] = 16'h7a7c;
initial mem[305] = 16'h7a41;
initial mem[306] = 16'h7a04;
initial mem[307] = 16'h79c7;
initial mem[308] = 16'h7989;
initial mem[309] = 16'h7949;
initial mem[310] = 16'h7908;
initial mem[311] = 16'h78c6;
initial mem[312] = 16'h7883;
initial mem[313] = 16'h783f;
initial mem[314] = 16'h77f9;
initial mem[315] = 16'h77b3;
initial mem[316] = 16'h776b;
initial mem[317] = 16'h7722;
initial mem[318] = 16'h76d8;
initial mem[319] = 16'h768d;
initial mem[320] = 16'h7640;
initial mem[321] = 16'h75f3;
initial mem[322] = 16'h75a4;
initial mem[323] = 16'h7554;
initial mem[324] = 16'h7503;
initial mem[325] = 16'h74b1;
initial mem[326] = 16'h745e;
initial mem[327] = 16'h740a;
initial mem[328] = 16'h73b5;
initial mem[329] = 16'h735e;
initial mem[330] = 16'h7306;
initial mem[331] = 16'h72ae;
initial mem[332] = 16'h7254;
initial mem[333] = 16'h71f9;
initial mem[334] = 16'h719d;
initial mem[335] = 16'h7140;
initial mem[336] = 16'h70e1;
initial mem[337] = 16'h7082;
initial mem[338] = 16'h7022;
initial mem[339] = 16'h6fc0;
initial mem[340] = 16'h6f5e;
initial mem[341] = 16'h6efa;
initial mem[342] = 16'h6e95;
initial mem[343] = 16'h6e30;
initial mem[344] = 16'h6dc9;
initial mem[345] = 16'h6d61;
initial mem[346] = 16'h6cf8;
initial mem[347] = 16'h6c8e;
initial mem[348] = 16'h6c23;
initial mem[349] = 16'h6bb7;
initial mem[350] = 16'h6b4a;
initial mem[351] = 16'h6adb;
initial mem[352] = 16'h6a6c;
initial mem[353] = 16'h69fc;
initial mem[354] = 16'h698b;
initial mem[355] = 16'h6919;
initial mem[356] = 16'h68a5;
initial mem[357] = 16'h6831;
initial mem[358] = 16'h67bc;
initial mem[359] = 16'h6745;
initial mem[360] = 16'h66ce;
initial mem[361] = 16'h6656;
initial mem[362] = 16'h65dd;
initial mem[363] = 16'h6562;
initial mem[364] = 16'h64e7;
initial mem[365] = 16'h646b;
initial mem[366] = 16'h63ee;
initial mem[367] = 16'h6370;
initial mem[368] = 16'h62f1;
initial mem[369] = 16'h6271;
initial mem[370] = 16'h61f0;
initial mem[371] = 16'h616e;
initial mem[372] = 16'h60eb;
initial mem[373] = 16'h6067;
initial mem[374] = 16'h5fe2;
initial mem[375] = 16'h5f5d;
initial mem[376] = 16'h5ed6;
initial mem[377] = 16'h5e4f;
initial mem[378] = 16'h5dc6;
initial mem[379] = 16'h5d3d;
initial mem[380] = 16'h5cb3;
initial mem[381] = 16'h5c28;
initial mem[382] = 16'h5b9c;
initial mem[383] = 16'h5b0f;
initial mem[384] = 16'h5a81;
initial mem[385] = 16'h59f3;
initial mem[386] = 16'h5963;
initial mem[387] = 16'h58d3;
initial mem[388] = 16'h5842;
initial mem[389] = 16'h57b0;
initial mem[390] = 16'h571d;
initial mem[391] = 16'h5689;
initial mem[392] = 16'h55f4;
initial mem[393] = 16'h555f;
initial mem[394] = 16'h54c9;
initial mem[395] = 16'h5432;
initial mem[396] = 16'h539a;
initial mem[397] = 16'h5301;
initial mem[398] = 16'h5268;
initial mem[399] = 16'h51ce;
initial mem[400] = 16'h5133;
initial mem[401] = 16'h5097;
initial mem[402] = 16'h4ffa;
initial mem[403] = 16'h4f5d;
initial mem[404] = 16'h4ebf;
initial mem[405] = 16'h4e20;
initial mem[406] = 16'h4d80;
initial mem[407] = 16'h4ce0;
initial mem[408] = 16'h4c3f;
initial mem[409] = 16'h4b9d;
initial mem[410] = 16'h4afa;
initial mem[411] = 16'h4a57;
initial mem[412] = 16'h49b3;
initial mem[413] = 16'h490e;
initial mem[414] = 16'h4869;
initial mem[415] = 16'h47c3;
initial mem[416] = 16'h471c;
initial mem[417] = 16'h4674;
initial mem[418] = 16'h45cc;
initial mem[419] = 16'h4523;
initial mem[420] = 16'h447a;
initial mem[421] = 16'h43d0;
initial mem[422] = 16'h4325;
initial mem[423] = 16'h4279;
initial mem[424] = 16'h41cd;
initial mem[425] = 16'h4120;
initial mem[426] = 16'h4073;
initial mem[427] = 16'h3fc5;
initial mem[428] = 16'h3f16;
initial mem[429] = 16'h3e67;
initial mem[430] = 16'h3db7;
initial mem[431] = 16'h3d07;
initial mem[432] = 16'h3c56;
initial mem[433] = 16'h3ba4;
initial mem[434] = 16'h3af2;
initial mem[435] = 16'h3a3f;
initial mem[436] = 16'h398c;
initial mem[437] = 16'h38d8;
initial mem[438] = 16'h3824;
initial mem[439] = 16'h376f;
initial mem[440] = 16'h36b9;
initial mem[441] = 16'h3603;
initial mem[442] = 16'h354d;
initial mem[443] = 16'h3496;
initial mem[444] = 16'h33de;
initial mem[445] = 16'h3326;
initial mem[446] = 16'h326d;
initial mem[447] = 16'h31b4;
initial mem[448] = 16'h30fb;
initial mem[449] = 16'h3041;
initial mem[450] = 16'h2f86;
initial mem[451] = 16'h2ecc;
initial mem[452] = 16'h2e10;
initial mem[453] = 16'h2d54;
initial mem[454] = 16'h2c98;
initial mem[455] = 16'h2bdb;
initial mem[456] = 16'h2b1e;
initial mem[457] = 16'h2a61;
initial mem[458] = 16'h29a3;
initial mem[459] = 16'h28e5;
initial mem[460] = 16'h2826;
initial mem[461] = 16'h2767;
initial mem[462] = 16'h26a7;
initial mem[463] = 16'h25e7;
initial mem[464] = 16'h2527;
initial mem[465] = 16'h2467;
initial mem[466] = 16'h23a6;
initial mem[467] = 16'h22e4;
initial mem[468] = 16'h2223;
initial mem[469] = 16'h2161;
initial mem[470] = 16'h209f;
initial mem[471] = 16'h1fdc;
initial mem[472] = 16'h1f19;
initial mem[473] = 16'h1e56;
initial mem[474] = 16'h1d93;
initial mem[475] = 16'h1ccf;
initial mem[476] = 16'h1c0b;
initial mem[477] = 16'h1b46;
initial mem[478] = 16'h1a82;
initial mem[479] = 16'h19bd;
initial mem[480] = 16'h18f8;
initial mem[481] = 16'h1833;
initial mem[482] = 16'h176d;
initial mem[483] = 16'h16a7;
initial mem[484] = 16'h15e1;
initial mem[485] = 16'h151b;
initial mem[486] = 16'h1455;
initial mem[487] = 16'h138e;
initial mem[488] = 16'h12c7;
initial mem[489] = 16'h1200;
initial mem[490] = 16'h1139;
initial mem[491] = 16'h1072;
initial mem[492] = 16'hfab;
initial mem[493] = 16'hee3;
initial mem[494] = 16'he1b;
initial mem[495] = 16'hd53;
initial mem[496] = 16'hc8b;
initial mem[497] = 16'hbc3;
initial mem[498] = 16'hafb;
initial mem[499] = 16'ha32;
initial mem[500] = 16'h96a;
initial mem[501] = 16'h8a1;
initial mem[502] = 16'h7d9;
initial mem[503] = 16'h710;
initial mem[504] = 16'h647;
initial mem[505] = 16'h57e;
initial mem[506] = 16'h4b6;
initial mem[507] = 16'h3ed;
initial mem[508] = 16'h324;
initial mem[509] = 16'h25b;
initial mem[510] = 16'h192;
initial mem[511] = 16'hc9;
initial mem[512] = 16'h0;
initial mem[513] = 16'hff37;
initial mem[514] = 16'hfe6e;
initial mem[515] = 16'hfda5;
initial mem[516] = 16'hfcdc;
initial mem[517] = 16'hfc13;
initial mem[518] = 16'hfb4a;
initial mem[519] = 16'hfa82;
initial mem[520] = 16'hf9b9;
initial mem[521] = 16'hf8f0;
initial mem[522] = 16'hf827;
initial mem[523] = 16'hf75f;
initial mem[524] = 16'hf696;
initial mem[525] = 16'hf5ce;
initial mem[526] = 16'hf505;
initial mem[527] = 16'hf43d;
initial mem[528] = 16'hf375;
initial mem[529] = 16'hf2ad;
initial mem[530] = 16'hf1e5;
initial mem[531] = 16'hf11d;
initial mem[532] = 16'hf055;
initial mem[533] = 16'hef8e;
initial mem[534] = 16'heec7;
initial mem[535] = 16'hee00;
initial mem[536] = 16'hed39;
initial mem[537] = 16'hec72;
initial mem[538] = 16'hebab;
initial mem[539] = 16'heae5;
initial mem[540] = 16'hea1f;
initial mem[541] = 16'he959;
initial mem[542] = 16'he893;
initial mem[543] = 16'he7cd;
initial mem[544] = 16'he708;
initial mem[545] = 16'he643;
initial mem[546] = 16'he57e;
initial mem[547] = 16'he4ba;
initial mem[548] = 16'he3f5;
initial mem[549] = 16'he331;
initial mem[550] = 16'he26d;
initial mem[551] = 16'he1aa;
initial mem[552] = 16'he0e7;
initial mem[553] = 16'he024;
initial mem[554] = 16'hdf61;
initial mem[555] = 16'hde9f;
initial mem[556] = 16'hdddd;
initial mem[557] = 16'hdd1c;
initial mem[558] = 16'hdc5a;
initial mem[559] = 16'hdb99;
initial mem[560] = 16'hdad9;
initial mem[561] = 16'hda19;
initial mem[562] = 16'hd959;
initial mem[563] = 16'hd899;
initial mem[564] = 16'hd7da;
initial mem[565] = 16'hd71b;
initial mem[566] = 16'hd65d;
initial mem[567] = 16'hd59f;
initial mem[568] = 16'hd4e2;
initial mem[569] = 16'hd425;
initial mem[570] = 16'hd368;
initial mem[571] = 16'hd2ac;
initial mem[572] = 16'hd1f0;
initial mem[573] = 16'hd134;
initial mem[574] = 16'hd07a;
initial mem[575] = 16'hcfbf;
initial mem[576] = 16'hcf05;
initial mem[577] = 16'hce4c;
initial mem[578] = 16'hcd93;
initial mem[579] = 16'hccda;
initial mem[580] = 16'hcc22;
initial mem[581] = 16'hcb6a;
initial mem[582] = 16'hcab3;
initial mem[583] = 16'hc9fd;
initial mem[584] = 16'hc947;
initial mem[585] = 16'hc891;
initial mem[586] = 16'hc7dc;
initial mem[587] = 16'hc728;
initial mem[588] = 16'hc674;
initial mem[589] = 16'hc5c1;
initial mem[590] = 16'hc50e;
initial mem[591] = 16'hc45c;
initial mem[592] = 16'hc3aa;
initial mem[593] = 16'hc2f9;
initial mem[594] = 16'hc249;
initial mem[595] = 16'hc199;
initial mem[596] = 16'hc0ea;
initial mem[597] = 16'hc03b;
initial mem[598] = 16'hbf8d;
initial mem[599] = 16'hbee0;
initial mem[600] = 16'hbe33;
initial mem[601] = 16'hbd87;
initial mem[602] = 16'hbcdb;
initial mem[603] = 16'hbc30;
initial mem[604] = 16'hbb86;
initial mem[605] = 16'hbadd;
initial mem[606] = 16'hba34;
initial mem[607] = 16'hb98c;
initial mem[608] = 16'hb8e4;
initial mem[609] = 16'hb83d;
initial mem[610] = 16'hb797;
initial mem[611] = 16'hb6f2;
initial mem[612] = 16'hb64d;
initial mem[613] = 16'hb5a9;
initial mem[614] = 16'hb506;
initial mem[615] = 16'hb463;
initial mem[616] = 16'hb3c1;
initial mem[617] = 16'hb320;
initial mem[618] = 16'hb280;
initial mem[619] = 16'hb1e0;
initial mem[620] = 16'hb141;
initial mem[621] = 16'hb0a3;
initial mem[622] = 16'hb006;
initial mem[623] = 16'haf69;
initial mem[624] = 16'haecd;
initial mem[625] = 16'hae32;
initial mem[626] = 16'had98;
initial mem[627] = 16'hacff;
initial mem[628] = 16'hac66;
initial mem[629] = 16'habce;
initial mem[630] = 16'hab37;
initial mem[631] = 16'haaa1;
initial mem[632] = 16'haa0c;
initial mem[633] = 16'ha977;
initial mem[634] = 16'ha8e3;
initial mem[635] = 16'ha850;
initial mem[636] = 16'ha7be;
initial mem[637] = 16'ha72d;
initial mem[638] = 16'ha69d;
initial mem[639] = 16'ha60d;
initial mem[640] = 16'ha57f;
initial mem[641] = 16'ha4f1;
initial mem[642] = 16'ha464;
initial mem[643] = 16'ha3d8;
initial mem[644] = 16'ha34d;
initial mem[645] = 16'ha2c3;
initial mem[646] = 16'ha23a;
initial mem[647] = 16'ha1b1;
initial mem[648] = 16'ha12a;
initial mem[649] = 16'ha0a3;
initial mem[650] = 16'ha01e;
initial mem[651] = 16'h9f99;
initial mem[652] = 16'h9f15;
initial mem[653] = 16'h9e92;
initial mem[654] = 16'h9e10;
initial mem[655] = 16'h9d8f;
initial mem[656] = 16'h9d0f;
initial mem[657] = 16'h9c90;
initial mem[658] = 16'h9c12;
initial mem[659] = 16'h9b95;
initial mem[660] = 16'h9b19;
initial mem[661] = 16'h9a9e;
initial mem[662] = 16'h9a23;
initial mem[663] = 16'h99aa;
initial mem[664] = 16'h9932;
initial mem[665] = 16'h98bb;
initial mem[666] = 16'h9844;
initial mem[667] = 16'h97cf;
initial mem[668] = 16'h975b;
initial mem[669] = 16'h96e7;
initial mem[670] = 16'h9675;
initial mem[671] = 16'h9604;
initial mem[672] = 16'h9594;
initial mem[673] = 16'h9525;
initial mem[674] = 16'h94b6;
initial mem[675] = 16'h9449;
initial mem[676] = 16'h93dd;
initial mem[677] = 16'h9372;
initial mem[678] = 16'h9308;
initial mem[679] = 16'h929f;
initial mem[680] = 16'h9237;
initial mem[681] = 16'h91d0;
initial mem[682] = 16'h916b;
initial mem[683] = 16'h9106;
initial mem[684] = 16'h90a2;
initial mem[685] = 16'h9040;
initial mem[686] = 16'h8fde;
initial mem[687] = 16'h8f7e;
initial mem[688] = 16'h8f1f;
initial mem[689] = 16'h8ec0;
initial mem[690] = 16'h8e63;
initial mem[691] = 16'h8e07;
initial mem[692] = 16'h8dac;
initial mem[693] = 16'h8d52;
initial mem[694] = 16'h8cfa;
initial mem[695] = 16'h8ca2;
initial mem[696] = 16'h8c4b;
initial mem[697] = 16'h8bf6;
initial mem[698] = 16'h8ba2;
initial mem[699] = 16'h8b4f;
initial mem[700] = 16'h8afd;
initial mem[701] = 16'h8aac;
initial mem[702] = 16'h8a5c;
initial mem[703] = 16'h8a0d;
initial mem[704] = 16'h89c0;
initial mem[705] = 16'h8973;
initial mem[706] = 16'h8928;
initial mem[707] = 16'h88de;
initial mem[708] = 16'h8895;
initial mem[709] = 16'h884d;
initial mem[710] = 16'h8807;
initial mem[711] = 16'h87c1;
initial mem[712] = 16'h877d;
initial mem[713] = 16'h873a;
initial mem[714] = 16'h86f8;
initial mem[715] = 16'h86b7;
initial mem[716] = 16'h8677;
initial mem[717] = 16'h8639;
initial mem[718] = 16'h85fc;
initial mem[719] = 16'h85bf;
initial mem[720] = 16'h8584;
initial mem[721] = 16'h854b;
initial mem[722] = 16'h8512;
initial mem[723] = 16'h84db;
initial mem[724] = 16'h84a4;
initial mem[725] = 16'h846f;
initial mem[726] = 16'h843c;
initial mem[727] = 16'h8409;
initial mem[728] = 16'h83d7;
initial mem[729] = 16'h83a7;
initial mem[730] = 16'h8378;
initial mem[731] = 16'h834a;
initial mem[732] = 16'h831e;
initial mem[733] = 16'h82f2;
initial mem[734] = 16'h82c8;
initial mem[735] = 16'h829f;
initial mem[736] = 16'h8277;
initial mem[737] = 16'h8250;
initial mem[738] = 16'h822b;
initial mem[739] = 16'h8207;
initial mem[740] = 16'h81e4;
initial mem[741] = 16'h81c2;
initial mem[742] = 16'h81a2;
initial mem[743] = 16'h8182;
initial mem[744] = 16'h8164;
initial mem[745] = 16'h8147;
initial mem[746] = 16'h812c;
initial mem[747] = 16'h8111;
initial mem[748] = 16'h80f8;
initial mem[749] = 16'h80e0;
initial mem[750] = 16'h80c9;
initial mem[751] = 16'h80b4;
initial mem[752] = 16'h809f;
initial mem[753] = 16'h808c;
initial mem[754] = 16'h807a;
initial mem[755] = 16'h806a;
initial mem[756] = 16'h805a;
initial mem[757] = 16'h804c;
initial mem[758] = 16'h803f;
initial mem[759] = 16'h8033;
initial mem[760] = 16'h8029;
initial mem[761] = 16'h8020;
initial mem[762] = 16'h8018;
initial mem[763] = 16'h8011;
initial mem[764] = 16'h800b;
initial mem[765] = 16'h8007;
initial mem[766] = 16'h8004;
initial mem[767] = 16'h8002;
initial mem[768] = 16'h8001;
initial mem[769] = 16'h8002;
initial mem[770] = 16'h8004;
initial mem[771] = 16'h8007;
initial mem[772] = 16'h800b;
initial mem[773] = 16'h8011;
initial mem[774] = 16'h8018;
initial mem[775] = 16'h8020;
initial mem[776] = 16'h8029;
initial mem[777] = 16'h8033;
initial mem[778] = 16'h803f;
initial mem[779] = 16'h804c;
initial mem[780] = 16'h805a;
initial mem[781] = 16'h806a;
initial mem[782] = 16'h807a;
initial mem[783] = 16'h808c;
initial mem[784] = 16'h809f;
initial mem[785] = 16'h80b4;
initial mem[786] = 16'h80c9;
initial mem[787] = 16'h80e0;
initial mem[788] = 16'h80f8;
initial mem[789] = 16'h8111;
initial mem[790] = 16'h812c;
initial mem[791] = 16'h8147;
initial mem[792] = 16'h8164;
initial mem[793] = 16'h8182;
initial mem[794] = 16'h81a2;
initial mem[795] = 16'h81c2;
initial mem[796] = 16'h81e4;
initial mem[797] = 16'h8207;
initial mem[798] = 16'h822b;
initial mem[799] = 16'h8250;
initial mem[800] = 16'h8277;
initial mem[801] = 16'h829f;
initial mem[802] = 16'h82c8;
initial mem[803] = 16'h82f2;
initial mem[804] = 16'h831e;
initial mem[805] = 16'h834a;
initial mem[806] = 16'h8378;
initial mem[807] = 16'h83a7;
initial mem[808] = 16'h83d7;
initial mem[809] = 16'h8409;
initial mem[810] = 16'h843c;
initial mem[811] = 16'h846f;
initial mem[812] = 16'h84a4;
initial mem[813] = 16'h84db;
initial mem[814] = 16'h8512;
initial mem[815] = 16'h854b;
initial mem[816] = 16'h8584;
initial mem[817] = 16'h85bf;
initial mem[818] = 16'h85fc;
initial mem[819] = 16'h8639;
initial mem[820] = 16'h8677;
initial mem[821] = 16'h86b7;
initial mem[822] = 16'h86f8;
initial mem[823] = 16'h873a;
initial mem[824] = 16'h877d;
initial mem[825] = 16'h87c1;
initial mem[826] = 16'h8807;
initial mem[827] = 16'h884d;
initial mem[828] = 16'h8895;
initial mem[829] = 16'h88de;
initial mem[830] = 16'h8928;
initial mem[831] = 16'h8973;
initial mem[832] = 16'h89c0;
initial mem[833] = 16'h8a0d;
initial mem[834] = 16'h8a5c;
initial mem[835] = 16'h8aac;
initial mem[836] = 16'h8afd;
initial mem[837] = 16'h8b4f;
initial mem[838] = 16'h8ba2;
initial mem[839] = 16'h8bf6;
initial mem[840] = 16'h8c4b;
initial mem[841] = 16'h8ca2;
initial mem[842] = 16'h8cfa;
initial mem[843] = 16'h8d52;
initial mem[844] = 16'h8dac;
initial mem[845] = 16'h8e07;
initial mem[846] = 16'h8e63;
initial mem[847] = 16'h8ec0;
initial mem[848] = 16'h8f1f;
initial mem[849] = 16'h8f7e;
initial mem[850] = 16'h8fde;
initial mem[851] = 16'h9040;
initial mem[852] = 16'h90a2;
initial mem[853] = 16'h9106;
initial mem[854] = 16'h916b;
initial mem[855] = 16'h91d0;
initial mem[856] = 16'h9237;
initial mem[857] = 16'h929f;
initial mem[858] = 16'h9308;
initial mem[859] = 16'h9372;
initial mem[860] = 16'h93dd;
initial mem[861] = 16'h9449;
initial mem[862] = 16'h94b6;
initial mem[863] = 16'h9525;
initial mem[864] = 16'h9594;
initial mem[865] = 16'h9604;
initial mem[866] = 16'h9675;
initial mem[867] = 16'h96e7;
initial mem[868] = 16'h975b;
initial mem[869] = 16'h97cf;
initial mem[870] = 16'h9844;
initial mem[871] = 16'h98bb;
initial mem[872] = 16'h9932;
initial mem[873] = 16'h99aa;
initial mem[874] = 16'h9a23;
initial mem[875] = 16'h9a9e;
initial mem[876] = 16'h9b19;
initial mem[877] = 16'h9b95;
initial mem[878] = 16'h9c12;
initial mem[879] = 16'h9c90;
initial mem[880] = 16'h9d0f;
initial mem[881] = 16'h9d8f;
initial mem[882] = 16'h9e10;
initial mem[883] = 16'h9e92;
initial mem[884] = 16'h9f15;
initial mem[885] = 16'h9f99;
initial mem[886] = 16'ha01e;
initial mem[887] = 16'ha0a3;
initial mem[888] = 16'ha12a;
initial mem[889] = 16'ha1b1;
initial mem[890] = 16'ha23a;
initial mem[891] = 16'ha2c3;
initial mem[892] = 16'ha34d;
initial mem[893] = 16'ha3d8;
initial mem[894] = 16'ha464;
initial mem[895] = 16'ha4f1;
initial mem[896] = 16'ha57f;
initial mem[897] = 16'ha60d;
initial mem[898] = 16'ha69d;
initial mem[899] = 16'ha72d;
initial mem[900] = 16'ha7be;
initial mem[901] = 16'ha850;
initial mem[902] = 16'ha8e3;
initial mem[903] = 16'ha977;
initial mem[904] = 16'haa0c;
initial mem[905] = 16'haaa1;
initial mem[906] = 16'hab37;
initial mem[907] = 16'habce;
initial mem[908] = 16'hac66;
initial mem[909] = 16'hacff;
initial mem[910] = 16'had98;
initial mem[911] = 16'hae32;
initial mem[912] = 16'haecd;
initial mem[913] = 16'haf69;
initial mem[914] = 16'hb006;
initial mem[915] = 16'hb0a3;
initial mem[916] = 16'hb141;
initial mem[917] = 16'hb1e0;
initial mem[918] = 16'hb280;
initial mem[919] = 16'hb320;
initial mem[920] = 16'hb3c1;
initial mem[921] = 16'hb463;
initial mem[922] = 16'hb506;
initial mem[923] = 16'hb5a9;
initial mem[924] = 16'hb64d;
initial mem[925] = 16'hb6f2;
initial mem[926] = 16'hb797;
initial mem[927] = 16'hb83d;
initial mem[928] = 16'hb8e4;
initial mem[929] = 16'hb98c;
initial mem[930] = 16'hba34;
initial mem[931] = 16'hbadd;
initial mem[932] = 16'hbb86;
initial mem[933] = 16'hbc30;
initial mem[934] = 16'hbcdb;
initial mem[935] = 16'hbd87;
initial mem[936] = 16'hbe33;
initial mem[937] = 16'hbee0;
initial mem[938] = 16'hbf8d;
initial mem[939] = 16'hc03b;
initial mem[940] = 16'hc0ea;
initial mem[941] = 16'hc199;
initial mem[942] = 16'hc249;
initial mem[943] = 16'hc2f9;
initial mem[944] = 16'hc3aa;
initial mem[945] = 16'hc45c;
initial mem[946] = 16'hc50e;
initial mem[947] = 16'hc5c1;
initial mem[948] = 16'hc674;
initial mem[949] = 16'hc728;
initial mem[950] = 16'hc7dc;
initial mem[951] = 16'hc891;
initial mem[952] = 16'hc947;
initial mem[953] = 16'hc9fd;
initial mem[954] = 16'hcab3;
initial mem[955] = 16'hcb6a;
initial mem[956] = 16'hcc22;
initial mem[957] = 16'hccda;
initial mem[958] = 16'hcd93;
initial mem[959] = 16'hce4c;
initial mem[960] = 16'hcf05;
initial mem[961] = 16'hcfbf;
initial mem[962] = 16'hd07a;
initial mem[963] = 16'hd134;
initial mem[964] = 16'hd1f0;
initial mem[965] = 16'hd2ac;
initial mem[966] = 16'hd368;
initial mem[967] = 16'hd425;
initial mem[968] = 16'hd4e2;
initial mem[969] = 16'hd59f;
initial mem[970] = 16'hd65d;
initial mem[971] = 16'hd71b;
initial mem[972] = 16'hd7da;
initial mem[973] = 16'hd899;
initial mem[974] = 16'hd959;
initial mem[975] = 16'hda19;
initial mem[976] = 16'hdad9;
initial mem[977] = 16'hdb99;
initial mem[978] = 16'hdc5a;
initial mem[979] = 16'hdd1c;
initial mem[980] = 16'hdddd;
initial mem[981] = 16'hde9f;
initial mem[982] = 16'hdf61;
initial mem[983] = 16'he024;
initial mem[984] = 16'he0e7;
initial mem[985] = 16'he1aa;
initial mem[986] = 16'he26d;
initial mem[987] = 16'he331;
initial mem[988] = 16'he3f5;
initial mem[989] = 16'he4ba;
initial mem[990] = 16'he57e;
initial mem[991] = 16'he643;
initial mem[992] = 16'he708;
initial mem[993] = 16'he7cd;
initial mem[994] = 16'he893;
initial mem[995] = 16'he959;
initial mem[996] = 16'hea1f;
initial mem[997] = 16'heae5;
initial mem[998] = 16'hebab;
initial mem[999] = 16'hec72;
initial mem[1000] = 16'hed39;
initial mem[1001] = 16'hee00;
initial mem[1002] = 16'heec7;
initial mem[1003] = 16'hef8e;
initial mem[1004] = 16'hf055;
initial mem[1005] = 16'hf11d;
initial mem[1006] = 16'hf1e5;
initial mem[1007] = 16'hf2ad;
initial mem[1008] = 16'hf375;
initial mem[1009] = 16'hf43d;
initial mem[1010] = 16'hf505;
initial mem[1011] = 16'hf5ce;
initial mem[1012] = 16'hf696;
initial mem[1013] = 16'hf75f;
initial mem[1014] = 16'hf827;
initial mem[1015] = 16'hf8f0;
initial mem[1016] = 16'hf9b9;
initial mem[1017] = 16'hfa82;
initial mem[1018] = 16'hfb4a;
initial mem[1019] = 16'hfc13;
initial mem[1020] = 16'hfcdc;
initial mem[1021] = 16'hfda5;
initial mem[1022] = 16'hfe6e;
initial mem[1023] = 16'hff37;
always @(posedge clk) begin
	data <= mem[addr];
end
endmodule

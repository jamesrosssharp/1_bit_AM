module noiseTable(input clk, input [9:0] addr, output reg [15:0] data);
reg [15:0] mem [0:1023];
initial mem[0] = 16'h1745;
initial mem[1] = 16'h12f8;
initial mem[2] = 16'h5d2;
initial mem[3] = 16'h196e;
initial mem[4] = 16'h146a;
initial mem[5] = 16'h1a09;
initial mem[6] = 16'hf409;
initial mem[7] = 16'h1651;
initial mem[8] = 16'he008;
initial mem[9] = 16'hec7;
initial mem[10] = 16'he958;
initial mem[11] = 16'heb1f;
initial mem[12] = 16'hefa4;
initial mem[13] = 16'hf629;
initial mem[14] = 16'h1c5e;
initial mem[15] = 16'h13d0;
initial mem[16] = 16'hf9c9;
initial mem[17] = 16'h1004;
initial mem[18] = 16'he7ad;
initial mem[19] = 16'he877;
initial mem[20] = 16'he39f;
initial mem[21] = 16'he43b;
initial mem[22] = 16'hff53;
initial mem[23] = 16'h2d8;
initial mem[24] = 16'he664;
initial mem[25] = 16'he391;
initial mem[26] = 16'h14da;
initial mem[27] = 16'h959;
initial mem[28] = 16'he4dc;
initial mem[29] = 16'h742;
initial mem[30] = 16'h17bd;
initial mem[31] = 16'hf8fd;
initial mem[32] = 16'hc57;
initial mem[33] = 16'hf2fe;
initial mem[34] = 16'hfc91;
initial mem[35] = 16'h15f4;
initial mem[36] = 16'hfe35;
initial mem[37] = 16'h17c0;
initial mem[38] = 16'h374;
initial mem[39] = 16'hd2d;
initial mem[40] = 16'hf95d;
initial mem[41] = 16'hea8b;
initial mem[42] = 16'hf80c;
initial mem[43] = 16'h46f;
initial mem[44] = 16'h5cd;
initial mem[45] = 16'h1a04;
initial mem[46] = 16'heee6;
initial mem[47] = 16'hf957;
initial mem[48] = 16'h1050;
initial mem[49] = 16'h1702;
initial mem[50] = 16'he640;
initial mem[51] = 16'hecb7;
initial mem[52] = 16'hf6c9;
initial mem[53] = 16'he68a;
initial mem[54] = 16'h1ceb;
initial mem[55] = 16'h1729;
initial mem[56] = 16'hf396;
initial mem[57] = 16'hf587;
initial mem[58] = 16'he578;
initial mem[59] = 16'h1e1;
initial mem[60] = 16'hfa57;
initial mem[61] = 16'h8fd;
initial mem[62] = 16'h4fe;
initial mem[63] = 16'h815;
initial mem[64] = 16'hbdb;
initial mem[65] = 16'hffab;
initial mem[66] = 16'he827;
initial mem[67] = 16'hf884;
initial mem[68] = 16'hfd5e;
initial mem[69] = 16'hb3b;
initial mem[70] = 16'h1399;
initial mem[71] = 16'h773;
initial mem[72] = 16'hc37;
initial mem[73] = 16'h1ae;
initial mem[74] = 16'he601;
initial mem[75] = 16'he322;
initial mem[76] = 16'he4af;
initial mem[77] = 16'hfa0;
initial mem[78] = 16'hf5b8;
initial mem[79] = 16'hf8aa;
initial mem[80] = 16'h5d7;
initial mem[81] = 16'hf448;
initial mem[82] = 16'he8b7;
initial mem[83] = 16'hf44b;
initial mem[84] = 16'hf2e6;
initial mem[85] = 16'hf814;
initial mem[86] = 16'h36e;
initial mem[87] = 16'hf58f;
initial mem[88] = 16'h6df;
initial mem[89] = 16'hedf0;
initial mem[90] = 16'h1e7d;
initial mem[91] = 16'hf03c;
initial mem[92] = 16'hf26a;
initial mem[93] = 16'hfb4;
initial mem[94] = 16'hfa3a;
initial mem[95] = 16'hc96;
initial mem[96] = 16'he8a1;
initial mem[97] = 16'hfad3;
initial mem[98] = 16'h4d1;
initial mem[99] = 16'he0e8;
initial mem[100] = 16'h1ca8;
initial mem[101] = 16'h28b;
initial mem[102] = 16'h71e;
initial mem[103] = 16'h1a06;
initial mem[104] = 16'h2d0;
initial mem[105] = 16'hf69b;
initial mem[106] = 16'hd82;
initial mem[107] = 16'h15e2;
initial mem[108] = 16'hfa61;
initial mem[109] = 16'he38b;
initial mem[110] = 16'h1bfe;
initial mem[111] = 16'h1fba;
initial mem[112] = 16'h786;
initial mem[113] = 16'hf50f;
initial mem[114] = 16'h1b93;
initial mem[115] = 16'he32f;
initial mem[116] = 16'h115a;
initial mem[117] = 16'hef43;
initial mem[118] = 16'hf704;
initial mem[119] = 16'h1eb;
initial mem[120] = 16'h134f;
initial mem[121] = 16'he859;
initial mem[122] = 16'hee14;
initial mem[123] = 16'he615;
initial mem[124] = 16'h140d;
initial mem[125] = 16'h6cc;
initial mem[126] = 16'h1391;
initial mem[127] = 16'h54d;
initial mem[128] = 16'h184b;
initial mem[129] = 16'hee03;
initial mem[130] = 16'hea24;
initial mem[131] = 16'h34f;
initial mem[132] = 16'h1628;
initial mem[133] = 16'h160c;
initial mem[134] = 16'hf3f3;
initial mem[135] = 16'hfc71;
initial mem[136] = 16'he9c9;
initial mem[137] = 16'h2c7;
initial mem[138] = 16'he36c;
initial mem[139] = 16'hfae2;
initial mem[140] = 16'he2f3;
initial mem[141] = 16'hffaa;
initial mem[142] = 16'h963;
initial mem[143] = 16'hf522;
initial mem[144] = 16'ha2f;
initial mem[145] = 16'hffd2;
initial mem[146] = 16'hf91c;
initial mem[147] = 16'hf9d6;
initial mem[148] = 16'hfa30;
initial mem[149] = 16'h31a;
initial mem[150] = 16'hff4;
initial mem[151] = 16'h384;
initial mem[152] = 16'hfcb0;
initial mem[153] = 16'hd6;
initial mem[154] = 16'h647;
initial mem[155] = 16'hf371;
initial mem[156] = 16'h4c5;
initial mem[157] = 16'hf3c2;
initial mem[158] = 16'h1e46;
initial mem[159] = 16'hf69d;
initial mem[160] = 16'he102;
initial mem[161] = 16'ha28;
initial mem[162] = 16'hf2fe;
initial mem[163] = 16'hff63;
initial mem[164] = 16'hf41e;
initial mem[165] = 16'hf345;
initial mem[166] = 16'hb4b;
initial mem[167] = 16'hf00a;
initial mem[168] = 16'hfeaf;
initial mem[169] = 16'hf799;
initial mem[170] = 16'he14c;
initial mem[171] = 16'h1093;
initial mem[172] = 16'h1fbf;
initial mem[173] = 16'hee14;
initial mem[174] = 16'hfbbb;
initial mem[175] = 16'he460;
initial mem[176] = 16'hf46b;
initial mem[177] = 16'he438;
initial mem[178] = 16'h1266;
initial mem[179] = 16'h1eba;
initial mem[180] = 16'h1a8c;
initial mem[181] = 16'h53b;
initial mem[182] = 16'h1c42;
initial mem[183] = 16'h1d1e;
initial mem[184] = 16'hcbd;
initial mem[185] = 16'h14b9;
initial mem[186] = 16'hec66;
initial mem[187] = 16'he363;
initial mem[188] = 16'h4ea;
initial mem[189] = 16'h426;
initial mem[190] = 16'he7b9;
initial mem[191] = 16'hc01;
initial mem[192] = 16'h15fc;
initial mem[193] = 16'hf923;
initial mem[194] = 16'hfde0;
initial mem[195] = 16'he24e;
initial mem[196] = 16'hf615;
initial mem[197] = 16'hfeee;
initial mem[198] = 16'he444;
initial mem[199] = 16'hfb7c;
initial mem[200] = 16'hfa91;
initial mem[201] = 16'h1593;
initial mem[202] = 16'h1b9f;
initial mem[203] = 16'h127e;
initial mem[204] = 16'hf125;
initial mem[205] = 16'hf2c;
initial mem[206] = 16'h1445;
initial mem[207] = 16'hef10;
initial mem[208] = 16'hf6c7;
initial mem[209] = 16'hf6d2;
initial mem[210] = 16'he185;
initial mem[211] = 16'he83c;
initial mem[212] = 16'he89f;
initial mem[213] = 16'h1b0;
initial mem[214] = 16'hf6ad;
initial mem[215] = 16'h8cd;
initial mem[216] = 16'he6a4;
initial mem[217] = 16'hd54;
initial mem[218] = 16'h1dd6;
initial mem[219] = 16'hd21;
initial mem[220] = 16'h137d;
initial mem[221] = 16'he79f;
initial mem[222] = 16'ha54;
initial mem[223] = 16'hf08e;
initial mem[224] = 16'he68;
initial mem[225] = 16'h1e40;
initial mem[226] = 16'heb4d;
initial mem[227] = 16'h1052;
initial mem[228] = 16'hfe10;
initial mem[229] = 16'hb29;
initial mem[230] = 16'h8dc;
initial mem[231] = 16'hf42d;
initial mem[232] = 16'hf31d;
initial mem[233] = 16'he353;
initial mem[234] = 16'hfdd1;
initial mem[235] = 16'haaf;
initial mem[236] = 16'h16c0;
initial mem[237] = 16'he0cc;
initial mem[238] = 16'h623;
initial mem[239] = 16'hff3;
initial mem[240] = 16'hebef;
initial mem[241] = 16'hff64;
initial mem[242] = 16'he01e;
initial mem[243] = 16'h13ca;
initial mem[244] = 16'h16e2;
initial mem[245] = 16'h4c4;
initial mem[246] = 16'he45;
initial mem[247] = 16'hf3e;
initial mem[248] = 16'he41c;
initial mem[249] = 16'h1a3;
initial mem[250] = 16'h166a;
initial mem[251] = 16'he1de;
initial mem[252] = 16'hed18;
initial mem[253] = 16'h1ce;
initial mem[254] = 16'he6c6;
initial mem[255] = 16'he16e;
initial mem[256] = 16'heb03;
initial mem[257] = 16'he3db;
initial mem[258] = 16'hbca;
initial mem[259] = 16'h96e;
initial mem[260] = 16'h2dc;
initial mem[261] = 16'hf4f5;
initial mem[262] = 16'hf054;
initial mem[263] = 16'h480;
initial mem[264] = 16'heb89;
initial mem[265] = 16'h1c6e;
initial mem[266] = 16'hf391;
initial mem[267] = 16'ha5;
initial mem[268] = 16'hf248;
initial mem[269] = 16'hef7e;
initial mem[270] = 16'h14b6;
initial mem[271] = 16'h1e25;
initial mem[272] = 16'hfead;
initial mem[273] = 16'he1df;
initial mem[274] = 16'hfb1a;
initial mem[275] = 16'hae5;
initial mem[276] = 16'h673;
initial mem[277] = 16'hfcaf;
initial mem[278] = 16'h17c1;
initial mem[279] = 16'h1aad;
initial mem[280] = 16'he61a;
initial mem[281] = 16'h5f8;
initial mem[282] = 16'h143a;
initial mem[283] = 16'he5a;
initial mem[284] = 16'he5f2;
initial mem[285] = 16'heeca;
initial mem[286] = 16'hf132;
initial mem[287] = 16'ha57;
initial mem[288] = 16'hf8b3;
initial mem[289] = 16'h4d3;
initial mem[290] = 16'he0ff;
initial mem[291] = 16'h1621;
initial mem[292] = 16'he087;
initial mem[293] = 16'hcc0;
initial mem[294] = 16'h1f9f;
initial mem[295] = 16'h1240;
initial mem[296] = 16'h1fe;
initial mem[297] = 16'h16f9;
initial mem[298] = 16'hf58e;
initial mem[299] = 16'he672;
initial mem[300] = 16'hffbc;
initial mem[301] = 16'hf6a6;
initial mem[302] = 16'h1cfc;
initial mem[303] = 16'hf73e;
initial mem[304] = 16'hfcf4;
initial mem[305] = 16'hf61a;
initial mem[306] = 16'h1aef;
initial mem[307] = 16'hf888;
initial mem[308] = 16'ha74;
initial mem[309] = 16'h1f71;
initial mem[310] = 16'hf4e5;
initial mem[311] = 16'h13f;
initial mem[312] = 16'h9fd;
initial mem[313] = 16'hf6f8;
initial mem[314] = 16'h187e;
initial mem[315] = 16'hadf;
initial mem[316] = 16'hfae7;
initial mem[317] = 16'h11ef;
initial mem[318] = 16'h1a7f;
initial mem[319] = 16'h14a9;
initial mem[320] = 16'hf60f;
initial mem[321] = 16'he226;
initial mem[322] = 16'hed18;
initial mem[323] = 16'hf3b8;
initial mem[324] = 16'hf0a3;
initial mem[325] = 16'hf71a;
initial mem[326] = 16'h116;
initial mem[327] = 16'h1ca4;
initial mem[328] = 16'he028;
initial mem[329] = 16'hf1a2;
initial mem[330] = 16'hef77;
initial mem[331] = 16'h1f52;
initial mem[332] = 16'h1dd6;
initial mem[333] = 16'h698;
initial mem[334] = 16'hced;
initial mem[335] = 16'he264;
initial mem[336] = 16'hfca8;
initial mem[337] = 16'hefc3;
initial mem[338] = 16'h1825;
initial mem[339] = 16'hf9ed;
initial mem[340] = 16'hea3a;
initial mem[341] = 16'hf93c;
initial mem[342] = 16'hf8f6;
initial mem[343] = 16'h1298;
initial mem[344] = 16'hfaac;
initial mem[345] = 16'hf373;
initial mem[346] = 16'h1029;
initial mem[347] = 16'h1126;
initial mem[348] = 16'h11c6;
initial mem[349] = 16'he1e1;
initial mem[350] = 16'he447;
initial mem[351] = 16'h1924;
initial mem[352] = 16'heda0;
initial mem[353] = 16'hea9a;
initial mem[354] = 16'h1909;
initial mem[355] = 16'he86e;
initial mem[356] = 16'ha1c;
initial mem[357] = 16'hed0d;
initial mem[358] = 16'hb63;
initial mem[359] = 16'h1258;
initial mem[360] = 16'h7cd;
initial mem[361] = 16'h1437;
initial mem[362] = 16'h4d0;
initial mem[363] = 16'h13dc;
initial mem[364] = 16'hfd28;
initial mem[365] = 16'hf240;
initial mem[366] = 16'he0a2;
initial mem[367] = 16'h68f;
initial mem[368] = 16'h19e8;
initial mem[369] = 16'h13ac;
initial mem[370] = 16'he71c;
initial mem[371] = 16'hfaa6;
initial mem[372] = 16'hd77;
initial mem[373] = 16'hf2ac;
initial mem[374] = 16'h171f;
initial mem[375] = 16'hfb9f;
initial mem[376] = 16'hfca0;
initial mem[377] = 16'he5ad;
initial mem[378] = 16'hec44;
initial mem[379] = 16'hebe4;
initial mem[380] = 16'h1222;
initial mem[381] = 16'h1f91;
initial mem[382] = 16'hef9e;
initial mem[383] = 16'hea0b;
initial mem[384] = 16'hfa24;
initial mem[385] = 16'he4c7;
initial mem[386] = 16'hf296;
initial mem[387] = 16'hd72;
initial mem[388] = 16'he112;
initial mem[389] = 16'he3ec;
initial mem[390] = 16'he43a;
initial mem[391] = 16'h710;
initial mem[392] = 16'hfa8c;
initial mem[393] = 16'h942;
initial mem[394] = 16'h37d;
initial mem[395] = 16'hee2;
initial mem[396] = 16'he7b7;
initial mem[397] = 16'h1ff5;
initial mem[398] = 16'hf205;
initial mem[399] = 16'hbbb;
initial mem[400] = 16'hb83;
initial mem[401] = 16'h1767;
initial mem[402] = 16'hebae;
initial mem[403] = 16'hf45d;
initial mem[404] = 16'hf452;
initial mem[405] = 16'hb0c;
initial mem[406] = 16'heb84;
initial mem[407] = 16'h3c1;
initial mem[408] = 16'ha6c;
initial mem[409] = 16'hf949;
initial mem[410] = 16'hee4a;
initial mem[411] = 16'hee12;
initial mem[412] = 16'h7c5;
initial mem[413] = 16'he956;
initial mem[414] = 16'he680;
initial mem[415] = 16'h1df4;
initial mem[416] = 16'hf9a8;
initial mem[417] = 16'h9ee;
initial mem[418] = 16'he167;
initial mem[419] = 16'he62c;
initial mem[420] = 16'h3ed;
initial mem[421] = 16'he9a3;
initial mem[422] = 16'hf7e9;
initial mem[423] = 16'he35d;
initial mem[424] = 16'hfc8f;
initial mem[425] = 16'he1b9;
initial mem[426] = 16'h1b7f;
initial mem[427] = 16'h705;
initial mem[428] = 16'hfd73;
initial mem[429] = 16'hfeb6;
initial mem[430] = 16'he0b;
initial mem[431] = 16'hffc4;
initial mem[432] = 16'he4d8;
initial mem[433] = 16'hc2a;
initial mem[434] = 16'h1597;
initial mem[435] = 16'hefd7;
initial mem[436] = 16'heb82;
initial mem[437] = 16'h1197;
initial mem[438] = 16'heb68;
initial mem[439] = 16'hfea8;
initial mem[440] = 16'h7d2;
initial mem[441] = 16'hf8e8;
initial mem[442] = 16'h3e4;
initial mem[443] = 16'hfafc;
initial mem[444] = 16'hf07c;
initial mem[445] = 16'hc6f;
initial mem[446] = 16'hff71;
initial mem[447] = 16'h175c;
initial mem[448] = 16'hfae9;
initial mem[449] = 16'he63d;
initial mem[450] = 16'h1d15;
initial mem[451] = 16'he76;
initial mem[452] = 16'h1ab5;
initial mem[453] = 16'he857;
initial mem[454] = 16'hfeda;
initial mem[455] = 16'h107;
initial mem[456] = 16'hee37;
initial mem[457] = 16'heee4;
initial mem[458] = 16'hee50;
initial mem[459] = 16'h15d0;
initial mem[460] = 16'hf646;
initial mem[461] = 16'hf593;
initial mem[462] = 16'hbfd;
initial mem[463] = 16'hfddd;
initial mem[464] = 16'h13ea;
initial mem[465] = 16'hf348;
initial mem[466] = 16'hef5e;
initial mem[467] = 16'h1599;
initial mem[468] = 16'h718;
initial mem[469] = 16'hf57a;
initial mem[470] = 16'hec07;
initial mem[471] = 16'h183f;
initial mem[472] = 16'hf5d9;
initial mem[473] = 16'hf93d;
initial mem[474] = 16'hf874;
initial mem[475] = 16'he09e;
initial mem[476] = 16'hf893;
initial mem[477] = 16'h1c7b;
initial mem[478] = 16'h1d2b;
initial mem[479] = 16'hf058;
initial mem[480] = 16'h1b8e;
initial mem[481] = 16'hfce0;
initial mem[482] = 16'hfe59;
initial mem[483] = 16'h477;
initial mem[484] = 16'h1746;
initial mem[485] = 16'hf8f0;
initial mem[486] = 16'hf1bd;
initial mem[487] = 16'h1310;
initial mem[488] = 16'h11a7;
initial mem[489] = 16'hfb05;
initial mem[490] = 16'hf3bf;
initial mem[491] = 16'h129;
initial mem[492] = 16'h132f;
initial mem[493] = 16'hf5cf;
initial mem[494] = 16'he6c2;
initial mem[495] = 16'h1b2f;
initial mem[496] = 16'h1999;
initial mem[497] = 16'hbff;
initial mem[498] = 16'h1aae;
initial mem[499] = 16'he231;
initial mem[500] = 16'h527;
initial mem[501] = 16'hf1b9;
initial mem[502] = 16'hba6;
initial mem[503] = 16'hfce5;
initial mem[504] = 16'hb64;
initial mem[505] = 16'hbd7;
initial mem[506] = 16'hf0b7;
initial mem[507] = 16'h174c;
initial mem[508] = 16'ha8f;
initial mem[509] = 16'hf3a7;
initial mem[510] = 16'he48;
initial mem[511] = 16'hfee4;
initial mem[512] = 16'he445;
initial mem[513] = 16'h1b67;
initial mem[514] = 16'hec0c;
initial mem[515] = 16'he2b3;
initial mem[516] = 16'he631;
initial mem[517] = 16'hed1a;
initial mem[518] = 16'h16af;
initial mem[519] = 16'heab2;
initial mem[520] = 16'h1a39;
initial mem[521] = 16'he8ba;
initial mem[522] = 16'h15c6;
initial mem[523] = 16'h1046;
initial mem[524] = 16'he7b8;
initial mem[525] = 16'heb50;
initial mem[526] = 16'h421;
initial mem[527] = 16'h5f0;
initial mem[528] = 16'hd56;
initial mem[529] = 16'h5de;
initial mem[530] = 16'hd57;
initial mem[531] = 16'h7aa;
initial mem[532] = 16'hf8e5;
initial mem[533] = 16'hf734;
initial mem[534] = 16'he614;
initial mem[535] = 16'hb3;
initial mem[536] = 16'hfc34;
initial mem[537] = 16'hedca;
initial mem[538] = 16'h18aa;
initial mem[539] = 16'hc89;
initial mem[540] = 16'ha10;
initial mem[541] = 16'he952;
initial mem[542] = 16'h159d;
initial mem[543] = 16'h1932;
initial mem[544] = 16'h7e4;
initial mem[545] = 16'hf698;
initial mem[546] = 16'hfd33;
initial mem[547] = 16'h58c;
initial mem[548] = 16'hedc4;
initial mem[549] = 16'hfbfd;
initial mem[550] = 16'heeb6;
initial mem[551] = 16'hf24;
initial mem[552] = 16'h1e1f;
initial mem[553] = 16'hf159;
initial mem[554] = 16'hea58;
initial mem[555] = 16'hbc4;
initial mem[556] = 16'he94a;
initial mem[557] = 16'h1f55;
initial mem[558] = 16'hf333;
initial mem[559] = 16'hed21;
initial mem[560] = 16'he2bc;
initial mem[561] = 16'he3e5;
initial mem[562] = 16'he965;
initial mem[563] = 16'hed08;
initial mem[564] = 16'hffbc;
initial mem[565] = 16'hf371;
initial mem[566] = 16'hed5d;
initial mem[567] = 16'h1f05;
initial mem[568] = 16'hf9d9;
initial mem[569] = 16'hf832;
initial mem[570] = 16'h1e8a;
initial mem[571] = 16'hfdc3;
initial mem[572] = 16'h831;
initial mem[573] = 16'hfac3;
initial mem[574] = 16'h18cb;
initial mem[575] = 16'h105e;
initial mem[576] = 16'h1519;
initial mem[577] = 16'h1634;
initial mem[578] = 16'h71d;
initial mem[579] = 16'hf8a7;
initial mem[580] = 16'h1e87;
initial mem[581] = 16'h2cd;
initial mem[582] = 16'heebe;
initial mem[583] = 16'hf158;
initial mem[584] = 16'he730;
initial mem[585] = 16'hf65f;
initial mem[586] = 16'heba7;
initial mem[587] = 16'he421;
initial mem[588] = 16'h1f9;
initial mem[589] = 16'h1cab;
initial mem[590] = 16'hdd3;
initial mem[591] = 16'hfb61;
initial mem[592] = 16'h12cc;
initial mem[593] = 16'he07c;
initial mem[594] = 16'he813;
initial mem[595] = 16'hebc9;
initial mem[596] = 16'hff9;
initial mem[597] = 16'h115;
initial mem[598] = 16'he8ef;
initial mem[599] = 16'he211;
initial mem[600] = 16'hf6b0;
initial mem[601] = 16'h16ec;
initial mem[602] = 16'h122d;
initial mem[603] = 16'hed8d;
initial mem[604] = 16'h17d2;
initial mem[605] = 16'hcac;
initial mem[606] = 16'he520;
initial mem[607] = 16'hf574;
initial mem[608] = 16'hbe0;
initial mem[609] = 16'hc81;
initial mem[610] = 16'hea67;
initial mem[611] = 16'h5db;
initial mem[612] = 16'hf37;
initial mem[613] = 16'h9f0;
initial mem[614] = 16'h1655;
initial mem[615] = 16'he114;
initial mem[616] = 16'he3ef;
initial mem[617] = 16'h1425;
initial mem[618] = 16'h362;
initial mem[619] = 16'he5bd;
initial mem[620] = 16'he578;
initial mem[621] = 16'hf32d;
initial mem[622] = 16'hf88a;
initial mem[623] = 16'hab;
initial mem[624] = 16'hebbd;
initial mem[625] = 16'hefa2;
initial mem[626] = 16'h11c9;
initial mem[627] = 16'heae6;
initial mem[628] = 16'hf547;
initial mem[629] = 16'hf5c9;
initial mem[630] = 16'he268;
initial mem[631] = 16'hff95;
initial mem[632] = 16'hf27c;
initial mem[633] = 16'hf9f3;
initial mem[634] = 16'h13bf;
initial mem[635] = 16'heb1a;
initial mem[636] = 16'h1cca;
initial mem[637] = 16'he993;
initial mem[638] = 16'h5d6;
initial mem[639] = 16'heba9;
initial mem[640] = 16'hecb;
initial mem[641] = 16'he44b;
initial mem[642] = 16'hfedd;
initial mem[643] = 16'he7a4;
initial mem[644] = 16'hf229;
initial mem[645] = 16'hf2ee;
initial mem[646] = 16'h43f;
initial mem[647] = 16'hf266;
initial mem[648] = 16'hfd59;
initial mem[649] = 16'hf39c;
initial mem[650] = 16'hea6c;
initial mem[651] = 16'h182d;
initial mem[652] = 16'hf939;
initial mem[653] = 16'h142b;
initial mem[654] = 16'he62;
initial mem[655] = 16'h12ea;
initial mem[656] = 16'hea16;
initial mem[657] = 16'he02c;
initial mem[658] = 16'he5e5;
initial mem[659] = 16'hf2cf;
initial mem[660] = 16'hec64;
initial mem[661] = 16'he530;
initial mem[662] = 16'hf214;
initial mem[663] = 16'he961;
initial mem[664] = 16'hef95;
initial mem[665] = 16'h8f;
initial mem[666] = 16'h828;
initial mem[667] = 16'hed40;
initial mem[668] = 16'hee10;
initial mem[669] = 16'hecd6;
initial mem[670] = 16'heaa8;
initial mem[671] = 16'hf730;
initial mem[672] = 16'h1e39;
initial mem[673] = 16'h1ae3;
initial mem[674] = 16'hd6f;
initial mem[675] = 16'hff5c;
initial mem[676] = 16'had6;
initial mem[677] = 16'h188;
initial mem[678] = 16'hf194;
initial mem[679] = 16'h17dc;
initial mem[680] = 16'hcff;
initial mem[681] = 16'h3f3;
initial mem[682] = 16'h1c96;
initial mem[683] = 16'h1e01;
initial mem[684] = 16'h173d;
initial mem[685] = 16'hfb97;
initial mem[686] = 16'h87e;
initial mem[687] = 16'he699;
initial mem[688] = 16'he2b1;
initial mem[689] = 16'hfd80;
initial mem[690] = 16'h16dc;
initial mem[691] = 16'h1c10;
initial mem[692] = 16'hd7e;
initial mem[693] = 16'hec1a;
initial mem[694] = 16'he911;
initial mem[695] = 16'he0cd;
initial mem[696] = 16'h1bac;
initial mem[697] = 16'hfb12;
initial mem[698] = 16'h1ba0;
initial mem[699] = 16'h5c0;
initial mem[700] = 16'hee98;
initial mem[701] = 16'he421;
initial mem[702] = 16'hfe7f;
initial mem[703] = 16'hf6a5;
initial mem[704] = 16'hf422;
initial mem[705] = 16'h14dd;
initial mem[706] = 16'hf077;
initial mem[707] = 16'h1e8c;
initial mem[708] = 16'hff2f;
initial mem[709] = 16'hfe04;
initial mem[710] = 16'h117c;
initial mem[711] = 16'h1fc4;
initial mem[712] = 16'hf551;
initial mem[713] = 16'he881;
initial mem[714] = 16'h10fc;
initial mem[715] = 16'he63b;
initial mem[716] = 16'hf1af;
initial mem[717] = 16'h1d6e;
initial mem[718] = 16'he3dd;
initial mem[719] = 16'hfb9b;
initial mem[720] = 16'hf561;
initial mem[721] = 16'he36a;
initial mem[722] = 16'hffd7;
initial mem[723] = 16'h58d;
initial mem[724] = 16'hf32e;
initial mem[725] = 16'hffc0;
initial mem[726] = 16'he55a;
initial mem[727] = 16'hf754;
initial mem[728] = 16'hf414;
initial mem[729] = 16'h1ca5;
initial mem[730] = 16'h173a;
initial mem[731] = 16'hee9a;
initial mem[732] = 16'he8f3;
initial mem[733] = 16'he0d1;
initial mem[734] = 16'h3c9;
initial mem[735] = 16'he365;
initial mem[736] = 16'he1ac;
initial mem[737] = 16'h44a;
initial mem[738] = 16'h189f;
initial mem[739] = 16'hfe44;
initial mem[740] = 16'h1ccc;
initial mem[741] = 16'h2d4;
initial mem[742] = 16'he81d;
initial mem[743] = 16'hc1d;
initial mem[744] = 16'h1c2c;
initial mem[745] = 16'he699;
initial mem[746] = 16'hf89d;
initial mem[747] = 16'he3f2;
initial mem[748] = 16'heef7;
initial mem[749] = 16'hfb5a;
initial mem[750] = 16'h1b7;
initial mem[751] = 16'hf43e;
initial mem[752] = 16'he0d6;
initial mem[753] = 16'he7a1;
initial mem[754] = 16'h469;
initial mem[755] = 16'hfdae;
initial mem[756] = 16'h134a;
initial mem[757] = 16'hf8cd;
initial mem[758] = 16'hfe25;
initial mem[759] = 16'h4b1;
initial mem[760] = 16'hf3aa;
initial mem[761] = 16'hed2f;
initial mem[762] = 16'hd1d;
initial mem[763] = 16'h90a;
initial mem[764] = 16'hf634;
initial mem[765] = 16'he119;
initial mem[766] = 16'h15fb;
initial mem[767] = 16'hf16;
initial mem[768] = 16'h1628;
initial mem[769] = 16'hef4;
initial mem[770] = 16'h8be;
initial mem[771] = 16'hf389;
initial mem[772] = 16'h1c30;
initial mem[773] = 16'h1b51;
initial mem[774] = 16'h223;
initial mem[775] = 16'h10c;
initial mem[776] = 16'hf414;
initial mem[777] = 16'hf1f9;
initial mem[778] = 16'h15b;
initial mem[779] = 16'hf690;
initial mem[780] = 16'hfece;
initial mem[781] = 16'he501;
initial mem[782] = 16'heee7;
initial mem[783] = 16'hf872;
initial mem[784] = 16'hfd97;
initial mem[785] = 16'he185;
initial mem[786] = 16'hf772;
initial mem[787] = 16'hfe91;
initial mem[788] = 16'hf1c2;
initial mem[789] = 16'hfd61;
initial mem[790] = 16'haf0;
initial mem[791] = 16'h197a;
initial mem[792] = 16'hfbc2;
initial mem[793] = 16'he474;
initial mem[794] = 16'he821;
initial mem[795] = 16'h1ced;
initial mem[796] = 16'hfd7f;
initial mem[797] = 16'hf1b9;
initial mem[798] = 16'heb89;
initial mem[799] = 16'hcb3;
initial mem[800] = 16'hf0a6;
initial mem[801] = 16'h177c;
initial mem[802] = 16'hf573;
initial mem[803] = 16'he6dc;
initial mem[804] = 16'hea07;
initial mem[805] = 16'hbb9;
initial mem[806] = 16'hf45c;
initial mem[807] = 16'hed56;
initial mem[808] = 16'haef;
initial mem[809] = 16'hfef4;
initial mem[810] = 16'h435;
initial mem[811] = 16'h6e5;
initial mem[812] = 16'h1a04;
initial mem[813] = 16'hea86;
initial mem[814] = 16'hfa1a;
initial mem[815] = 16'hf191;
initial mem[816] = 16'heb82;
initial mem[817] = 16'h1b50;
initial mem[818] = 16'hfc73;
initial mem[819] = 16'h1512;
initial mem[820] = 16'h187d;
initial mem[821] = 16'h1fdd;
initial mem[822] = 16'hf2ae;
initial mem[823] = 16'h9f8;
initial mem[824] = 16'hef2;
initial mem[825] = 16'h1ee5;
initial mem[826] = 16'hb0f;
initial mem[827] = 16'he7b5;
initial mem[828] = 16'h8ed;
initial mem[829] = 16'h59a;
initial mem[830] = 16'hf8d4;
initial mem[831] = 16'heaa2;
initial mem[832] = 16'he4c0;
initial mem[833] = 16'hed9d;
initial mem[834] = 16'hee7b;
initial mem[835] = 16'h911;
initial mem[836] = 16'he1dc;
initial mem[837] = 16'he788;
initial mem[838] = 16'he9f7;
initial mem[839] = 16'heb1d;
initial mem[840] = 16'hfbea;
initial mem[841] = 16'h1302;
initial mem[842] = 16'h101d;
initial mem[843] = 16'he801;
initial mem[844] = 16'hf87e;
initial mem[845] = 16'h1a0e;
initial mem[846] = 16'h10be;
initial mem[847] = 16'h17b3;
initial mem[848] = 16'hfd4e;
initial mem[849] = 16'hea2;
initial mem[850] = 16'h188a;
initial mem[851] = 16'hee4c;
initial mem[852] = 16'hf8fa;
initial mem[853] = 16'hf14e;
initial mem[854] = 16'h4c1;
initial mem[855] = 16'he5cd;
initial mem[856] = 16'hff75;
initial mem[857] = 16'hdf5;
initial mem[858] = 16'hf47;
initial mem[859] = 16'h193f;
initial mem[860] = 16'hd1;
initial mem[861] = 16'heb1e;
initial mem[862] = 16'he267;
initial mem[863] = 16'hf7e4;
initial mem[864] = 16'h639;
initial mem[865] = 16'h1f8a;
initial mem[866] = 16'h18c4;
initial mem[867] = 16'h1447;
initial mem[868] = 16'he08a;
initial mem[869] = 16'h117c;
initial mem[870] = 16'h3d7;
initial mem[871] = 16'hed87;
initial mem[872] = 16'hf4db;
initial mem[873] = 16'hfa29;
initial mem[874] = 16'hf895;
initial mem[875] = 16'hd6;
initial mem[876] = 16'hf590;
initial mem[877] = 16'h117c;
initial mem[878] = 16'h1b43;
initial mem[879] = 16'h1c6d;
initial mem[880] = 16'h1b9c;
initial mem[881] = 16'hfbed;
initial mem[882] = 16'hfcf;
initial mem[883] = 16'hf969;
initial mem[884] = 16'h1b3f;
initial mem[885] = 16'h1147;
initial mem[886] = 16'hfe40;
initial mem[887] = 16'h1b69;
initial mem[888] = 16'he5f3;
initial mem[889] = 16'hd94;
initial mem[890] = 16'h1873;
initial mem[891] = 16'h443;
initial mem[892] = 16'hefde;
initial mem[893] = 16'hf0c3;
initial mem[894] = 16'h1a06;
initial mem[895] = 16'h1ccd;
initial mem[896] = 16'he8e6;
initial mem[897] = 16'hfe23;
initial mem[898] = 16'h946;
initial mem[899] = 16'h102e;
initial mem[900] = 16'hf469;
initial mem[901] = 16'hf8f0;
initial mem[902] = 16'hec01;
initial mem[903] = 16'he85a;
initial mem[904] = 16'hf17b;
initial mem[905] = 16'hc2b;
initial mem[906] = 16'hfe3;
initial mem[907] = 16'h1bb2;
initial mem[908] = 16'he357;
initial mem[909] = 16'ha33;
initial mem[910] = 16'hffc5;
initial mem[911] = 16'h9ec;
initial mem[912] = 16'hc0a;
initial mem[913] = 16'h603;
initial mem[914] = 16'hebb4;
initial mem[915] = 16'heec2;
initial mem[916] = 16'hf3e5;
initial mem[917] = 16'hfef3;
initial mem[918] = 16'hfe2f;
initial mem[919] = 16'h98d;
initial mem[920] = 16'hfacd;
initial mem[921] = 16'hdd2;
initial mem[922] = 16'h1c89;
initial mem[923] = 16'hebba;
initial mem[924] = 16'hff63;
initial mem[925] = 16'h1f16;
initial mem[926] = 16'hfa5;
initial mem[927] = 16'h576;
initial mem[928] = 16'hef07;
initial mem[929] = 16'h8e5;
initial mem[930] = 16'hfea4;
initial mem[931] = 16'hf5d8;
initial mem[932] = 16'hf2a9;
initial mem[933] = 16'hea9;
initial mem[934] = 16'he99a;
initial mem[935] = 16'he264;
initial mem[936] = 16'hf283;
initial mem[937] = 16'h1b6d;
initial mem[938] = 16'hb53;
initial mem[939] = 16'h1c36;
initial mem[940] = 16'he39e;
initial mem[941] = 16'he123;
initial mem[942] = 16'h14bc;
initial mem[943] = 16'h1ab3;
initial mem[944] = 16'h6f9;
initial mem[945] = 16'he358;
initial mem[946] = 16'hf529;
initial mem[947] = 16'he094;
initial mem[948] = 16'h12d3;
initial mem[949] = 16'hf617;
initial mem[950] = 16'hfa67;
initial mem[951] = 16'hfd7a;
initial mem[952] = 16'he021;
initial mem[953] = 16'h1e10;
initial mem[954] = 16'hce8;
initial mem[955] = 16'hfbfa;
initial mem[956] = 16'hc77;
initial mem[957] = 16'h1a84;
initial mem[958] = 16'hfbaa;
initial mem[959] = 16'hea13;
initial mem[960] = 16'hdf4;
initial mem[961] = 16'he853;
initial mem[962] = 16'hf4b1;
initial mem[963] = 16'hf415;
initial mem[964] = 16'h1127;
initial mem[965] = 16'hf48a;
initial mem[966] = 16'h13fb;
initial mem[967] = 16'h1543;
initial mem[968] = 16'h130e;
initial mem[969] = 16'hef3b;
initial mem[970] = 16'h16f2;
initial mem[971] = 16'h1986;
initial mem[972] = 16'hf253;
initial mem[973] = 16'h8bf;
initial mem[974] = 16'h122;
initial mem[975] = 16'he1c8;
initial mem[976] = 16'hf893;
initial mem[977] = 16'he041;
initial mem[978] = 16'hb85;
initial mem[979] = 16'h1c1b;
initial mem[980] = 16'hf295;
initial mem[981] = 16'h12fa;
initial mem[982] = 16'h10e;
initial mem[983] = 16'hc7e;
initial mem[984] = 16'hf2d9;
initial mem[985] = 16'h1838;
initial mem[986] = 16'hf443;
initial mem[987] = 16'h1500;
initial mem[988] = 16'h90d;
initial mem[989] = 16'h730;
initial mem[990] = 16'h7f5;
initial mem[991] = 16'heda3;
initial mem[992] = 16'h90e;
initial mem[993] = 16'h25f;
initial mem[994] = 16'h198c;
initial mem[995] = 16'he6f8;
initial mem[996] = 16'heaa7;
initial mem[997] = 16'hf9ff;
initial mem[998] = 16'h1bd5;
initial mem[999] = 16'he46d;
initial mem[1000] = 16'hf7b9;
initial mem[1001] = 16'he554;
initial mem[1002] = 16'he0ec;
initial mem[1003] = 16'hef05;
initial mem[1004] = 16'heeac;
initial mem[1005] = 16'hf6eb;
initial mem[1006] = 16'he78;
initial mem[1007] = 16'h1ef9;
initial mem[1008] = 16'he2c9;
initial mem[1009] = 16'h1bad;
initial mem[1010] = 16'h1804;
initial mem[1011] = 16'h805;
initial mem[1012] = 16'he080;
initial mem[1013] = 16'he2fc;
initial mem[1014] = 16'haab;
initial mem[1015] = 16'hf008;
initial mem[1016] = 16'h1946;
initial mem[1017] = 16'h1d96;
initial mem[1018] = 16'h547;
initial mem[1019] = 16'hffc1;
initial mem[1020] = 16'he847;
initial mem[1021] = 16'he423;
initial mem[1022] = 16'h413;
initial mem[1023] = 16'h1b0d;
always @(posedge clk) begin
	data <= mem[addr];
end
endmodule
